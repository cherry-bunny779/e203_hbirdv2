`define RISCV_FORMAL
`define RISCV_FORMAL_NRET 1
`define RISCV_FORMAL_XLEN 32
`define RISCV_FORMAL_ILEN 32
`include "e203_defines.v"

module e203_hbirdv2 (
  // Preserve all original ports and macros from e203_cpu_top
  output [`E203_PC_SIZE-1:0] inspect_pc,
  output inspect_dbg_irq,
  output inspect_mem_cmd_valid,
  output inspect_mem_cmd_ready,
  output inspect_mem_rsp_valid,
  output inspect_mem_rsp_ready,
  output inspect_core_clk,
  output core_csr_clk,
  output core_wfi,
  output tm_stop,
  input  [`E203_PC_SIZE-1:0] pc_rtvec,
  output dbg_irq_r,
  output [`E203_PC_SIZE-1:0] cmt_dpc,
  output cmt_dpc_ena,
  output [2:0] cmt_dcause,
  output cmt_dcause_ena,
  output wr_dcsr_ena,
  output wr_dpc_ena,
  output wr_dscratch_ena,
  output [31:0] wr_csr_nxt,
  input  [31:0] dcsr_r,
  input  [`E203_PC_SIZE-1:0] dpc_r,
  input  [31:0] dscratch_r,
  input  dbg_mode,
  input  dbg_halt_r,
  input  dbg_step_r,
  input  dbg_ebreakm_r,
  input  dbg_stopcycle,
  input  dbg_irq_a,
  input  [`E203_HART_ID_W-1:0] core_mhartid,
  input  ext_irq_a,
  input  sft_irq_a,
  input  tmr_irq_a,
  input  tcm_sd,
  input  tcm_ds,
`ifdef E203_HAS_ITCM_EXTITF
  input  ext2itcm_icb_cmd_valid,
  output ext2itcm_icb_cmd_ready,
  input  [`E203_ITCM_ADDR_WIDTH-1:0] ext2itcm_icb_cmd_addr,
  input  ext2itcm_icb_cmd_read,
  input  [`E203_XLEN-1:0] ext2itcm_icb_cmd_wdata,
  input  [`E203_XLEN/8-1:0] ext2itcm_icb_cmd_wmask,
  output ext2itcm_icb_rsp_valid,
  input  ext2itcm_icb_rsp_ready,
  output ext2itcm_icb_rsp_err,
  output [`E203_XLEN-1:0] ext2itcm_icb_rsp_rdata,
`endif
`ifdef E203_HAS_DTCM_EXTITF
  input  ext2dtcm_icb_cmd_valid,
  output ext2dtcm_icb_cmd_ready,
  input  [`E203_DTCM_ADDR_WIDTH-1:0] ext2dtcm_icb_cmd_addr,
  input  ext2dtcm_icb_cmd_read,
  input  [`E203_XLEN-1:0] ext2dtcm_icb_cmd_wdata,
  input  [`E203_XLEN/8-1:0] ext2dtcm_icb_cmd_wmask,
  output ext2dtcm_icb_rsp_valid,
  input  ext2dtcm_icb_rsp_ready,
  output ext2dtcm_icb_rsp_err,
  output [`E203_XLEN-1:0] ext2dtcm_icb_rsp_rdata,
`endif
  output ppi_icb_cmd_valid,
  input  ppi_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0] ppi_icb_cmd_addr,
  output ppi_icb_cmd_read,
  output [`E203_XLEN-1:0] ppi_icb_cmd_wdata,
  output [`E203_XLEN/8-1:0] ppi_icb_cmd_wmask,
  input  ppi_icb_rsp_valid,
  output ppi_icb_rsp_ready,
  input  ppi_icb_rsp_err,
  input  [`E203_XLEN-1:0] ppi_icb_rsp_rdata,
  output clint_icb_cmd_valid,
  input  clint_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0] clint_icb_cmd_addr,
  output clint_icb_cmd_read,
  output [`E203_XLEN-1:0] clint_icb_cmd_wdata,
  output [`E203_XLEN/8-1:0] clint_icb_cmd_wmask,
  input  clint_icb_rsp_valid,
  output clint_icb_rsp_ready,
  input  clint_icb_rsp_err,
  input  [`E203_XLEN-1:0] clint_icb_rsp_rdata,
  output plic_icb_cmd_valid,
  input  plic_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0] plic_icb_cmd_addr,
  output plic_icb_cmd_read,
  output [`E203_XLEN-1:0] plic_icb_cmd_wdata,
  output [`E203_XLEN/8-1:0] plic_icb_cmd_wmask,
  input  plic_icb_rsp_valid,
  output plic_icb_rsp_ready,
  input  plic_icb_rsp_err,
  input  [`E203_XLEN-1:0] plic_icb_rsp_rdata,
  output fio_icb_cmd_valid,
  input  fio_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0] fio_icb_cmd_addr,
  output fio_icb_cmd_read,
  output [`E203_XLEN-1:0] fio_icb_cmd_wdata,
  output [`E203_XLEN/8-1:0] fio_icb_cmd_wmask,
  input  fio_icb_rsp_valid,
  output fio_icb_rsp_ready,
  input  fio_icb_rsp_err,
  input  [`E203_XLEN-1:0] fio_icb_rsp_rdata,
  output mem_icb_cmd_valid,
  input  mem_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0] mem_icb_cmd_addr,
  output mem_icb_cmd_read,
  output [`E203_XLEN-1:0] mem_icb_cmd_wdata,
  output [`E203_XLEN/8-1:0] mem_icb_cmd_wmask,
  input  mem_icb_rsp_valid,
  output mem_icb_rsp_ready,
  input  mem_icb_rsp_err,
  input  [`E203_XLEN-1:0] mem_icb_rsp_rdata,
  input  test_mode,
  input  clk,
  input  rst_n
);

e203_cpu_top u_e203_cpu_top(
  .inspect_pc(inspect_pc),
  .inspect_dbg_irq(inspect_dbg_irq),
  .inspect_mem_cmd_valid(inspect_mem_cmd_valid),
  .inspect_mem_cmd_ready(inspect_mem_cmd_ready),
  .inspect_mem_rsp_valid(inspect_mem_rsp_valid),
  .inspect_mem_rsp_ready(inspect_mem_rsp_ready),
  .inspect_core_clk(inspect_core_clk),
  .core_csr_clk(core_csr_clk),
  .core_wfi(core_wfi),
  .tm_stop(tm_stop),
  .pc_rtvec(pc_rtvec),
  .dbg_irq_r(dbg_irq_r),
  .cmt_dpc(cmt_dpc),
  .cmt_dpc_ena(cmt_dpc_ena),
  .cmt_dcause(cmt_dcause),
  .cmt_dcause_ena(cmt_dcause_ena),
  .wr_dcsr_ena(wr_dcsr_ena),
  .wr_dpc_ena(wr_dpc_ena),
  .wr_dscratch_ena(wr_dscratch_ena),
  .wr_csr_nxt(wr_csr_nxt),
  .dcsr_r(dcsr_r),
  .dpc_r(dpc_r),
  .dscratch_r(dscratch_r),
  .dbg_mode(dbg_mode),
  .dbg_halt_r(dbg_halt_r),
  .dbg_step_r(dbg_step_r),
  .dbg_ebreakm_r(dbg_ebreakm_r),
  .dbg_stopcycle(dbg_stopcycle),
  .dbg_irq_a(dbg_irq_a),
  .core_mhartid(core_mhartid),
  .ext_irq_a(ext_irq_a),
  .sft_irq_a(sft_irq_a),
  .tmr_irq_a(tmr_irq_a),
  .tcm_sd(tcm_sd),
  .tcm_ds(tcm_ds),
`ifdef E203_HAS_ITCM_EXTITF
  .ext2itcm_icb_cmd_valid(ext2itcm_icb_cmd_valid),
  .ext2itcm_icb_cmd_ready(ext2itcm_icb_cmd_ready),
  .ext2itcm_icb_cmd_addr(ext2itcm_icb_cmd_addr),
  .ext2itcm_icb_cmd_read(ext2itcm_icb_cmd_read),
  .ext2itcm_icb_cmd_wdata(ext2itcm_icb_cmd_wdata),
  .ext2itcm_icb_cmd_wmask(ext2itcm_icb_cmd_wmask),
  .ext2itcm_icb_rsp_valid(ext2itcm_icb_rsp_valid),
  .ext2itcm_icb_rsp_ready(ext2itcm_icb_rsp_ready),
  .ext2itcm_icb_rsp_err(ext2itcm_icb_rsp_err),
  .ext2itcm_icb_rsp_rdata(ext2itcm_icb_rsp_rdata),
`endif
`ifdef E203_HAS_DTCM_EXTITF
  .ext2dtcm_icb_cmd_valid(ext2dtcm_icb_cmd_valid),
  .ext2dtcm_icb_cmd_ready(ext2dtcm_icb_cmd_ready),
  .ext2dtcm_icb_cmd_addr(ext2dtcm_icb_cmd_addr),
  .ext2dtcm_icb_cmd_read(ext2dtcm_icb_cmd_read),
  .ext2dtcm_icb_cmd_wdata(ext2dtcm_icb_cmd_wdata),
  .ext2dtcm_icb_cmd_wmask(ext2dtcm_icb_cmd_wmask),
  .ext2dtcm_icb_rsp_valid(ext2dtcm_icb_rsp_valid),
  .ext2dtcm_icb_rsp_ready(ext2dtcm_icb_rsp_ready),
  .ext2dtcm_icb_rsp_err(ext2dtcm_icb_rsp_err),
  .ext2dtcm_icb_rsp_rdata(ext2dtcm_icb_rsp_rdata),
`endif
  .ppi_icb_cmd_valid(ppi_icb_cmd_valid),
  .ppi_icb_cmd_ready(ppi_icb_cmd_ready),
  .ppi_icb_cmd_addr(ppi_icb_cmd_addr),
  .ppi_icb_cmd_read(ppi_icb_cmd_read),
  .ppi_icb_cmd_wdata(ppi_icb_cmd_wdata),
  .ppi_icb_cmd_wmask(ppi_icb_cmd_wmask),
  .ppi_icb_rsp_valid(ppi_icb_rsp_valid),
  .ppi_icb_rsp_ready(ppi_icb_rsp_ready),
  .ppi_icb_rsp_err(ppi_icb_rsp_err),
  .ppi_icb_rsp_rdata(ppi_icb_rsp_rdata),
  .clint_icb_cmd_valid(clint_icb_cmd_valid),
  .clint_icb_cmd_ready(clint_icb_cmd_ready),
  .clint_icb_cmd_addr(clint_icb_cmd_addr),
  .clint_icb_cmd_read(clint_icb_cmd_read),
  .clint_icb_cmd_wdata(clint_icb_cmd_wdata),
  .clint_icb_cmd_wmask(clint_icb_cmd_wmask),
  .clint_icb_rsp_valid(clint_icb_rsp_valid),
  .clint_icb_rsp_ready(clint_icb_rsp_ready),
  .clint_icb_rsp_err(clint_icb_rsp_err),
  .clint_icb_rsp_rdata(clint_icb_rsp_rdata),
  .plic_icb_cmd_valid(plic_icb_cmd_valid),
  .plic_icb_cmd_ready(plic_icb_cmd_ready),
  .plic_icb_cmd_addr(plic_icb_cmd_addr),
  .plic_icb_cmd_read(plic_icb_cmd_read),
  .plic_icb_cmd_wdata(plic_icb_cmd_wdata),
  .plic_icb_cmd_wmask(plic_icb_cmd_wmask),
  .plic_icb_rsp_valid(plic_icb_rsp_valid),
  .plic_icb_rsp_ready(plic_icb_rsp_ready),
  .plic_icb_rsp_err(plic_icb_rsp_err),
  .plic_icb_rsp_rdata(plic_icb_rsp_rdata),
  .fio_icb_cmd_valid(fio_icb_cmd_valid),
  .fio_icb_cmd_ready(fio_icb_cmd_ready),
  .fio_icb_cmd_addr(fio_icb_cmd_addr),
  .fio_icb_cmd_read(fio_icb_cmd_read),
  .fio_icb_cmd_wdata(fio_icb_cmd_wdata),
  .fio_icb_cmd_wmask(fio_icb_cmd_wmask),
  .fio_icb_rsp_valid(fio_icb_rsp_valid),
  .fio_icb_rsp_ready(fio_icb_rsp_ready),
  .fio_icb_rsp_err(fio_icb_rsp_err),
  .fio_icb_rsp_rdata(fio_icb_rsp_rdata),
  .mem_icb_cmd_valid(mem_icb_cmd_valid),
  .mem_icb_cmd_ready(mem_icb_cmd_ready),
  .mem_icb_cmd_addr(mem_icb_cmd_addr),
  .mem_icb_cmd_read(mem_icb_cmd_read),
  .mem_icb_cmd_wdata(mem_icb_cmd_wdata),
  .mem_icb_cmd_wmask(mem_icb_cmd_wmask),
  .mem_icb_rsp_valid(mem_icb_rsp_valid),
  .mem_icb_rsp_ready(mem_icb_rsp_ready),
  .mem_icb_rsp_err(mem_icb_rsp_err),
  .mem_icb_rsp_rdata(mem_icb_rsp_rdata),
  .test_mode(test_mode),
  .clk(clk),
  .rst_n(rst_n)
);

endmodule