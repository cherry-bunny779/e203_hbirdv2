always @* if (!reset) cover (channel[0].cnt_insns == 2);

