`define RISCV_FORMAL
`define RISCV_FORMAL_NRET 1
`define RISCV_FORMAL_XLEN 32
`define RISCV_FORMAL_ILEN 32
`define RISCV_FORMAL_RESET_CYCLES 1
`define RISCV_FORMAL_CHECK_CYCLE 15
`define RISCV_FORMAL_CHANNEL_IDX 0
`define RISCV_FORMAL_CHECKER rvfi_insn_check
`define RISCV_FORMAL_INSN_MODEL rvfi_insn_c_j
`define RISCV_FORMAL_COMPRESSED
`define RISCV_FORMAL_ALIGNED_MEM
`define RISCV_FORMAL_ALTOPS
`define RISCV_FORMAL_UMODE
`define PICORV32_TESTBUG_NONE
`define DEBUGNETS
`include "rvfi_macros.vh"

